//"
//
//
//"
//"
`include "i2c_if.sv"
`include "i2c_transaction.sv"
`include "i2c_sequence.sv"
`include "i2c_sequencer.sv"
`include "i2c_driver.sv"
`include "i2c_monitor.sv"
`include "monitor2.sv"
`include "i2c_agent.sv"
`include "i2c_freq_sb.sv"
`include "i2c_env.sv"
`include "i2c_test.sv"
//"
